module FakePrefetch(
  input         clock,
  input         reset,
  output        pf_train_ready,
  input         pf_train_valid,
  input  [20:0] pf_train_bits_tag,
  input  [8:0]  pf_train_bits_set,
  input         pf_train_bits_needT,
  input  [6:0]  pf_train_bits_source,
  input         pf_req_ready,
  output        pf_req_valid,
  output [20:0] pf_req_bits_tag,
  output [8:0]  pf_req_bits_set,
  output        pf_req_bits_needT,
  output [6:0]  pf_req_bits_source,
  output        pf_req_bits_isBOP,
  output        pf_resp_ready,
  input         pf_resp_valid,
  input  [20:0] pf_resp_bits_tag,
  input  [8:0]  pf_resp_bits_set,
  input         pf_recv_addr_valid,
  input  [63:0] pf_recv_addr_bits,
  input         pf_l2_pf_en
);
  pf_SppPrefetch spp (
    .clock(clock),
    .reset(reset),
    .io_train_ready(pf_train_ready),
    .io_train_valid(pf_train_valid),
    .io_train_bits_tag(pf_train_bits_tag),
    .io_train_bits_set(pf_train_bits_set),
    .io_train_bits_needT(pf_train_bits_needT),
    .io_train_bits_source(pf_train_bits_source),
    .io_req_ready(pf_req_ready),
    .io_req_valid(pf_req_valid),
    .io_req_bits_tag(pf_req_bits_tag),
    .io_req_bits_set(pf_req_bits_set),
    .io_req_bits_needT(pf_req_bits_needT),
    .io_req_bits_source(pf_req_bits_source),
    .io_req_bits_isBOP(pf_req_bits_isBOP),
    .io_resp_ready(pf_resp_ready),
    .io_resp_valid(pf_reso_valid),
    .io_resp_bits_tag(pf_resp_bits_tag),
    .io_resp_bits_set(pf_resp_bits_set)
  );
endmodule